//////////////////////////////////////////////////////////////////////////////////
// Exercise #5 
// Student Name: Akshay Pal
// Date: 9th June 2020
//
//  Description: In this exercise, you need to implement a UK traffic lights 
//  sequencing system. 
//
//  inputs:
//           clk
//
//  outputs:
//           red, amber, green
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 100ps

module lights (
	input clk,
	output reg red,
	output reg amber,
	output reg green
	);

	



